module ST_DPHD_HIPERF_2048x32m4_Tlmr (ATP,CK1,CK2,CSN1,CSN2,IG1,IG2,INITN,MTCK,
 SCTRLI1,SCTRLI2,SCTRLO1,SCTRLO2,SDLI1,SDLI2,SDLO1,SDLO2,SDRI1,SDRI2,
 SDRO1,SDRO2,SE,STDBY1,STDBY2,TBIST,TBYPASS,TCSN1,TCSN2,TED1,
 TED2,TOD1,TOD2,TP,TWEN1,TWEN2,WEN1,WEN2,A1,A2,
 D1,D2,Q1,Q2,TA1,TA2 );
 input ATP,CK1,CK2,CSN1,CSN2,IG1,IG2,INITN,MTCK,
 SCTRLI1,SCTRLI2,SDLI1,SDLI2,SDRI1,SDRI2,SE,STDBY1,STDBY2,TBIST,
 TBYPASS,TCSN1,TCSN2,TED1,TED2,TOD1,TOD2,TP,TWEN1,TWEN2,
 WEN1,WEN2;
 input [10:0] A1;
 input [10:0] A2;
 input [31:0] D1;
 input [31:0] D2;
 input [10:0] TA1;
 input [10:0] TA2;
 output SCTRLO1,SCTRLO2,SDLO1,SDLO2,SDRO1,SDRO2;
 output [31:0] Q1;
 output [31:0] Q2;
endmodule
