module ST_SPHD_HIPERF_1024x32m4_Tlmr (ATP,CK,CSN,IG,INITN,SCTRLI,SCTRLO,SDLI,SDLO,
 SDRI,SDRO,SE,STDBY,TBIST,TBYPASS,TCSN,TED,TOD,TWEN,
 WEN,A,D,Q,TA );
 input ATP,CK,CSN,IG,INITN,SCTRLI,SDLI,SDRI,SE,
 STDBY,TBIST,TBYPASS,TCSN,TED,TOD,TWEN,WEN;
 input [9:0] A;
 input [31:0] D;
 input [9:0] TA;
 output SCTRLO,SDLO,SDRO;
 output [31:0] Q;
endmodule
module ST_SPHD_HIPERF_2048x32m8_Tlmr (ATP,CK,CSN,IG,INITN,SCTRLI,SCTRLO,SDLI,SDLO,
 SDRI,SDRO,SE,STDBY,TBIST,TBYPASS,TCSN,TED,TOD,TWEN,
 WEN,A,D,Q,TA );
 input ATP,CK,CSN,IG,INITN,SCTRLI,SDLI,SDRI,SE,
 STDBY,TBIST,TBYPASS,TCSN,TED,TOD,TWEN,WEN;
 input [10:0] A;
 input [31:0] D;
 input [10:0] TA;
 output SCTRLO,SDLO,SDRO;
 output [31:0] Q;
endmodule
module ST_SPHD_HIPERF_3072x32m8_Tlmr (ATP,CK,CSN,IG,INITN,SCTRLI,SCTRLO,SDLI,SDLO,
 SDRI,SDRO,SE,STDBY,TBIST,TBYPASS,TCSN,TED,TOD,TWEN,
 WEN,A,D,Q,TA );
 input ATP,CK,CSN,IG,INITN,SCTRLI,SDLI,SDRI,SE,
 STDBY,TBIST,TBYPASS,TCSN,TED,TOD,TWEN,WEN;
 input [11:0] A;
 input [31:0] D;
 input [11:0] TA;
 output SCTRLO,SDLO,SDRO;
 output [31:0] Q;
endmodule
module ST_SPHD_HIPERF_4096x32m8_Tlmr_HIPERF_CUT (ATP,CK,CSN,IG,INITN,SCTRLI,SCTRLO,SDLI,SDLO,
 SDRI,SDRO,SE,STDBY,TBIST,TBYPASS,TCSN,TED,TOD,TWEN,
 WEN,A,D,Q,TA );
 input ATP,CK,CSN,IG,INITN,SCTRLI,SDLI,SDRI,SE,
 STDBY,TBIST,TBYPASS,TCSN,TED,TOD,TWEN,WEN;
 input [11:0] A;
 input [31:0] D;
 input [11:0] TA;
 output SCTRLO,SDLO,SDRO;
 output [31:0] Q;
endmodule
